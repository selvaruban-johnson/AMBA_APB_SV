
`include "amba_packet.sv"
`include "amba_generator.sv"
`include "amba_driver.sv"
`include "intf.sv"
`include "amba_apb.v"
`include "Probe_Packet.sv"
`include "Probe_Intf.sv"
`include "amba_monitor.sv"
`include "amba_coverage.sv"
`include "amba_scoreboard.sv"
`include "amba_environment.sv"
`include "amba_test.sv"