class Probe_Packet;

		logic psel,penable,pwrite;
		logic [7 : 0] paddr,pwdata,prdata;
		logic pready;


	function void pre_randomize();
		
	endfunction

	function void post_randomize();
		
	endfunction

endclass